library verilog;
use verilog.vl_types.all;
entity Hackathon_vlg_vec_tst is
end Hackathon_vlg_vec_tst;
